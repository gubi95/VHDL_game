--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   17:01:15 04/15/2017
-- Design Name:   
-- Module Name:   C:/Users/Admin/Documents/VHDL_game/game/vgaTest.vhd
-- Project Name:  game
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: VGA
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY vgaTest IS
END vgaTest;
 
ARCHITECTURE behavior OF vgaTest IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT VGA
    PORT(
         Clk : IN  std_logic;
         RGB : IN  std_logic_vector(2 downto 0);
         R : OUT  std_logic;
         G : OUT  std_logic;
         B : OUT  std_logic;
         HS : OUT  std_logic;
         VS : OUT  std_logic;
         frameEnded : OUT  std_logic;
         runADC : OUT  std_logic;
         dac : OUT  std_logic_vector(7 downto 0);
         currXPos : OUT  std_logic_vector(9 downto 0);
         currYPos : OUT  std_logic_vector(9 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal Clk : std_logic := '0';
   signal RGB : std_logic_vector(2 downto 0) := (others => '0');

 	--Outputs
   signal R : std_logic;
   signal G : std_logic;
   signal B : std_logic;
   signal HS : std_logic;
   signal VS : std_logic;
   signal frameEnded : std_logic;
   signal runADC : std_logic;
   signal dac : std_logic_vector(7 downto 0);
   signal currXPos : std_logic_vector(9 downto 0);
   signal currYPos : std_logic_vector(9 downto 0);

   -- Clock period definitions
   constant Clk_period : time := 20 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: VGA PORT MAP (
          Clk => Clk,
          RGB => RGB,
          R => R,
          G => G,
          B => B,
          HS => HS,
          VS => VS,
          frameEnded => frameEnded,
          runADC => runADC,
          dac => dac,
          currXPos => currXPos,
          currYPos => currYPos
        );

   -- Clock process definitions
   Clk_process :process
   begin
		Clk <= '0';
		wait for Clk_period/2;
		Clk <= '1';
		wait for Clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for Clk_period*10;

      -- insert stimulus here
			RGB <= "111";

      wait;
   end process;

END;
